`timescale 1ns / 1ps

module layer_2#(
DATA_WIDTH = 32
)(
input logic [DATA_WIDTH-1:0] data0,   // 채널 0의 입력 데이터
    input logic [DATA_WIDTH-1:0] data1,   // 채널 1의 입력 데이터
    input logic [DATA_WIDTH-1:0] data2,   // 채널 2의 입력 데이터
    input logic [DATA_WIDTH-1:0] data3,   // 채널 3의 입력 데이터
    input logic [DATA_WIDTH-1:0] data4,   // 채널 4의 입력 데이터
    input logic [DATA_WIDTH-1:0] data5,   // 채널 5의 입력 데이터
    input logic [DATA_WIDTH-1:0] data6,   // 채널 6의 입력 데이터
    input logic [DATA_WIDTH-1:0] data7,   // 채널 7의 입력 데이터
    input logic [DATA_WIDTH-1:0] data8,   // 채널 8의 입력 데이터
    input logic [DATA_WIDTH-1:0] data9,   // 채널 9의 입력 데이터
    input logic [DATA_WIDTH-1:0] data10,  // 채널 10의 입력 데이터
    input logic [DATA_WIDTH-1:0] data11,  // 채널 11의 입력 데이터
    input logic [DATA_WIDTH-1:0] data12,  // 채널 12의 입력 데이터
    input logic [DATA_WIDTH-1:0] data13,  // 채널 13의 입력 데이터
    input logic [DATA_WIDTH-1:0] data14,  // 채널 14의 입력 데이터
    input logic [DATA_WIDTH-1:0] data15,  // 채널 15의 입력 데이터
    input logic [DATA_WIDTH-1:0] data16,  // 채널 16의 입력 데이터
    input logic [DATA_WIDTH-1:0] data17,  // 채널 17의 입력 데이터
    input logic [DATA_WIDTH-1:0] data18,  // 채널 18의 입력 데이터
    input logic [DATA_WIDTH-1:0] data19,  // 채널 19의 입력 데이터
    input logic [DATA_WIDTH-1:0] data20,  // 채널 20의 입력 데이터
    input logic [DATA_WIDTH-1:0] data21,  // 채널 21의 입력 데이터
    input logic [DATA_WIDTH-1:0] data22,  // 채널 22의 입력 데이터
    input logic [DATA_WIDTH-1:0] data23,  // 채널 23의 입력 데이터
    input logic [DATA_WIDTH-1:0] data24,  // 채널 24의 입력 데이터
    input logic [DATA_WIDTH-1:0] data25,  // 채널 25의 입력 데이터
    input logic [DATA_WIDTH-1:0] data26,  // 채널 26의 입력 데이터
    input logic [DATA_WIDTH-1:0] data27,  // 채널 27의 입력 데이터
    input logic [DATA_WIDTH-1:0] data28,  // 채널 28의 입력 데이터
    input logic [DATA_WIDTH-1:0] data29,  // 채널 29의 입력 데이터
    input logic [DATA_WIDTH-1:0] data30,  // 채널 30의 입력 데이터
    input logic [DATA_WIDTH-1:0] data31,
    input valid_in,
    input clk,
    input rst_n,
    output reg [31:0] data_out_1,
    output reg [31:0] data_out_2,
    output reg [31:0] data_out_3,
    output reg [31:0] data_out_4,
    output reg [31:0] data_out_5,
    output reg [31:0] data_out_6,
    output reg [31:0] data_out_7,
    output reg [31:0] data_out_8,
    output reg [31:0] data_out_9,
    output reg [31:0] data_out_10,
    output reg [31:0] data_out_11,
    output reg [31:0] data_out_12,
    output reg [31:0] data_out_13,
    output reg [31:0] data_out_14,
    output reg [31:0] data_out_15,
    output reg [31:0] data_out_16,
    output reg [31:0] data_out_17,
    output reg [31:0] data_out_18,
    output reg [31:0] data_out_19,
    output reg [31:0] data_out_20,
    output reg [31:0] data_out_21,
    output reg [31:0] data_out_22,
    output reg [31:0] data_out_23,
    output reg [31:0] data_out_24,
    output reg [31:0] data_out_25,
    output reg [31:0] data_out_26,
    output reg [31:0] data_out_27,
    output reg [31:0] data_out_28,
    output reg [31:0] data_out_29,
    output reg [31:0] data_out_30,
    output reg [31:0] data_out_31,
    output reg [31:0] data_out_32,
    output reg [31:0] data_out_33,
    output reg [31:0] data_out_34,
    output reg [31:0] data_out_35,
    output reg [31:0] data_out_36,
    output reg [31:0] data_out_37,
    output reg [31:0] data_out_38,
    output reg [31:0] data_out_39,
    output reg [31:0] data_out_40,
    output reg [31:0] data_out_41,
    output reg [31:0] data_out_42,
    output reg [31:0] data_out_43,
    output reg [31:0] data_out_44,
    output reg [31:0] data_out_45,
    output reg [31:0] data_out_46,
    output reg [31:0] data_out_47,
    output reg [31:0] data_out_48,
    output reg [31:0] data_out_49,
    output reg [31:0] data_out_50,
    output reg [31:0] data_out_51,
    output reg [31:0] data_out_52,
    output reg [31:0] data_out_53,
    output reg [31:0] data_out_54,
    output reg [31:0] data_out_55,
    output reg [31:0] data_out_56,
    output reg [31:0] data_out_57,
    output reg [31:0] data_out_58,
    output reg [31:0] data_out_59,
    output reg [31:0] data_out_60,
    output reg [31:0] data_out_61,
    output reg [31:0] data_out_62,
    output reg [31:0] data_out_63,
    output reg [31:0] data_out_64,      
    output reg valid_out_layer2
    
    );
    
    
reg valid_out_input_buffer;
 reg [31:0] buffer0 [0:16][0:12];  // 채널 0의 버퍼
    reg [31:0] buffer1 [0:16][0:12];  // 채널 1의 버퍼
    reg [31:0] buffer2 [0:16][0:12];  // 채널 2의 버퍼
    reg [31:0] buffer3 [0:16][0:12];  // 채널 3의 버퍼
    reg [31:0] buffer4 [0:16][0:12];  // 채널 4의 버퍼
    reg [31:0] buffer5 [0:16][0:12];  // 채널 5의 버퍼
    reg [31:0] buffer6 [0:16][0:12];  // 채널 6의 버퍼
    reg [31:0] buffer7 [0:16][0:12];  // 채널 7의 버퍼
    reg [31:0] buffer8 [0:16][0:12];  // 채널 8의 버퍼
    reg [31:0] buffer9 [0:16][0:12];  // 채널 9의 버퍼
    reg [31:0] buffer10 [0:16][0:12]; // 채널 10의 버퍼
    reg [31:0] buffer11 [0:16][0:12]; // 채널 11의 버퍼
    reg [31:0] buffer12 [0:16][0:12]; // 채널 12의 버퍼
    reg [31:0] buffer13 [0:16][0:12]; // 채널 13의 버퍼
    reg [31:0] buffer14 [0:16][0:12]; // 채널 14의 버퍼
    reg [31:0] buffer15 [0:16][0:12]; // 채널 15의 버퍼
    reg [31:0] buffer16 [0:16][0:12]; // 채널 16의 버퍼
    reg [31:0] buffer17 [0:16][0:12]; // 채널 17의 버퍼
    reg [31:0] buffer18 [0:16][0:12]; // 채널 18의 버퍼
    reg [31:0] buffer19 [0:16][0:12]; // 채널 19의 버퍼
    reg [31:0] buffer20 [0:16][0:12]; // 채널 20의 버퍼
    reg [31:0] buffer21 [0:16][0:12]; // 채널 21의 버퍼
    reg [31:0] buffer22 [0:16][0:12]; // 채널 22의 버퍼
    reg [31:0] buffer23 [0:16][0:12]; // 채널 23의 버퍼
    reg [31:0] buffer24 [0:16][0:12]; // 채널 24의 버퍼
    reg [31:0] buffer25 [0:16][0:12]; // 채널 25의 버퍼
    reg [31:0] buffer26 [0:16][0:12]; // 채널 26의 버퍼
    reg [31:0] buffer27 [0:16][0:12]; // 채널 27의 버퍼
    reg [31:0] buffer28 [0:16][0:12]; // 채널 28의 버퍼
    reg [31:0] buffer29 [0:16][0:12]; // 채널 29의 버퍼
    reg [31:0] buffer30 [0:16][0:12]; // 채널 30의 버퍼
    reg [31:0] buffer31 [0:16][0:12]; // 채널 31의 버퍼    
    
    reg valid_out_zero_padding_second;
    reg [31:0] padded0  [0:18][0:14];  // 패딩 0
    reg [31:0] padded1  [0:18][0:14];  // 패딩 1
    reg [31:0] padded2  [0:18][0:14];  // 패딩 2
    reg [31:0] padded3  [0:18][0:14];  // 패딩 3
    reg [31:0] padded4  [0:18][0:14];  // 패딩 4
    reg [31:0] padded5  [0:18][0:14];  // 패딩 5
    reg [31:0] padded6  [0:18][0:14];  // 패딩 6
    reg [31:0] padded7  [0:18][0:14];  // 패딩 7
    reg [31:0] padded8  [0:18][0:14];  // 패딩 8
    reg [31:0] padded9  [0:18][0:14];  // 패딩 9
    reg [31:0] padded10 [0:18][0:14];  // 패딩 10
    reg [31:0] padded11 [0:18][0:14];  // 패딩 11
    reg [31:0] padded12 [0:18][0:14];  // 패딩 12
    reg [31:0] padded13 [0:18][0:14];  // 패딩 13
    reg [31:0] padded14 [0:18][0:14];  // 패딩 14
    reg [31:0] padded15 [0:18][0:14];  // 패딩 15
    reg [31:0] padded16 [0:18][0:14];  // 패딩 16
    reg [31:0] padded17 [0:18][0:14];  // 패딩 17
    reg [31:0] padded18 [0:18][0:14];  // 패딩 18
    reg [31:0] padded19 [0:18][0:14];  // 패딩 19
    reg [31:0] padded20 [0:18][0:14];  // 패딩 20
    reg [31:0] padded21 [0:18][0:14];  // 패딩 21
    reg [31:0] padded22 [0:18][0:14];  // 패딩 22
    reg [31:0] padded23 [0:18][0:14];  // 패딩 23
    reg [31:0] padded24 [0:18][0:14];  // 패딩 24
    reg [31:0] padded25 [0:18][0:14];  // 패딩 25
    reg [31:0] padded26 [0:18][0:14];  // 패딩 26
    reg [31:0] padded27 [0:18][0:14];  // 패딩 27
    reg [31:0] padded28 [0:18][0:14];  // 패딩 28
    reg [31:0] padded29 [0:18][0:14];  // 패딩 29
    reg [31:0] padded30 [0:18][0:14];  // 패딩 30
    reg [31:0] padded31 [0:18][0:14];  // 패딩 31
    
    reg valid_out_threebythree;
    reg [DATA_WIDTH-1:0] patch [0:2][0:2];
    
    reg [31:0] data_out_conv2 [0:63];
    reg valid_out_conv2;
    
    reg [31:0] data_out_conv2_accum [0:63];
    reg valid_out_conv2_accum;
    
    reg [31:0] data_out_relu2 [0:63];
    reg valid_out_relu2;    
    
    reg [31:0] data_out_buf_1  [0:1][0:1];
reg [31:0] data_out_buf_2  [0:1][0:1];
reg [31:0] data_out_buf_3  [0:1][0:1];
reg [31:0] data_out_buf_4  [0:1][0:1];
reg [31:0] data_out_buf_5  [0:1][0:1];
reg [31:0] data_out_buf_6  [0:1][0:1];
reg [31:0] data_out_buf_7  [0:1][0:1];
reg [31:0] data_out_buf_8  [0:1][0:1];
reg [31:0] data_out_buf_9  [0:1][0:1];
reg [31:0] data_out_buf_10 [0:1][0:1];
reg [31:0] data_out_buf_11 [0:1][0:1];
reg [31:0] data_out_buf_12 [0:1][0:1];
reg [31:0] data_out_buf_13 [0:1][0:1];
reg [31:0] data_out_buf_14 [0:1][0:1];
reg [31:0] data_out_buf_15 [0:1][0:1];
reg [31:0] data_out_buf_16 [0:1][0:1];
reg [31:0] data_out_buf_17 [0:1][0:1];
reg [31:0] data_out_buf_18 [0:1][0:1];
reg [31:0] data_out_buf_19 [0:1][0:1];
reg [31:0] data_out_buf_20 [0:1][0:1];
reg [31:0] data_out_buf_21 [0:1][0:1];
reg [31:0] data_out_buf_22 [0:1][0:1];
reg [31:0] data_out_buf_23 [0:1][0:1];
reg [31:0] data_out_buf_24 [0:1][0:1];
reg [31:0] data_out_buf_25 [0:1][0:1];
reg [31:0] data_out_buf_26 [0:1][0:1];
reg [31:0] data_out_buf_27 [0:1][0:1];
reg [31:0] data_out_buf_28 [0:1][0:1];
reg [31:0] data_out_buf_29 [0:1][0:1];
reg [31:0] data_out_buf_30 [0:1][0:1];
reg [31:0] data_out_buf_31 [0:1][0:1];
reg [31:0] data_out_buf_32 [0:1][0:1];
reg [31:0] data_out_buf_33 [0:1][0:1];
reg [31:0] data_out_buf_34 [0:1][0:1];
reg [31:0] data_out_buf_35 [0:1][0:1];
reg [31:0] data_out_buf_36 [0:1][0:1];
reg [31:0] data_out_buf_37 [0:1][0:1];
reg [31:0] data_out_buf_38 [0:1][0:1];
reg [31:0] data_out_buf_39 [0:1][0:1];
reg [31:0] data_out_buf_40 [0:1][0:1];
reg [31:0] data_out_buf_41 [0:1][0:1];
reg [31:0] data_out_buf_42 [0:1][0:1];
reg [31:0] data_out_buf_43 [0:1][0:1];
reg [31:0] data_out_buf_44 [0:1][0:1];
reg [31:0] data_out_buf_45 [0:1][0:1];
reg [31:0] data_out_buf_46 [0:1][0:1];
reg [31:0] data_out_buf_47 [0:1][0:1];
reg [31:0] data_out_buf_48 [0:1][0:1];
reg [31:0] data_out_buf_49 [0:1][0:1];
reg [31:0] data_out_buf_50 [0:1][0:1];
reg [31:0] data_out_buf_51 [0:1][0:1];
reg [31:0] data_out_buf_52 [0:1][0:1];
reg [31:0] data_out_buf_53 [0:1][0:1];
reg [31:0] data_out_buf_54 [0:1][0:1];
reg [31:0] data_out_buf_55 [0:1][0:1];
reg [31:0] data_out_buf_56 [0:1][0:1];
reg [31:0] data_out_buf_57 [0:1][0:1];
reg [31:0] data_out_buf_58 [0:1][0:1];
reg [31:0] data_out_buf_59 [0:1][0:1];
reg [31:0] data_out_buf_60 [0:1][0:1];
reg [31:0] data_out_buf_61 [0:1][0:1];
reg [31:0] data_out_buf_62 [0:1][0:1];
reg [31:0] data_out_buf_63 [0:1][0:1];
reg [31:0] data_out_buf_64 [0:1][0:1];
reg valid_out_channel_buffer2;

input_buffer #(
.DATA_WIDTH(32),
.CHANNELS(32),
.WIDTH(13),
.HEIGHT(17)
)input_buffer(
.valid_in(valid_in),
.data0(data0),
.data1(data1),
.data2(data2),
.data3(data3),
.data4(data4),
.data5(data5),
.data6(data6),
.data7(data7),
.data8(data8),
.data9(data9),
.data10(data10),
.data11(data11),
.data12(data12),
.data13(data13),
.data14(data14),
.data15(data15),
.data16(data16),
.data17(data17),
.data18(data18),
.data19(data19),
.data20(data20),
.data21(data21),
.data22(data22),
.data23(data23),
.data24(data24),
.data25(data25),
.data26(data26),
.data27(data27),
.data28(data28),
.data29(data29),
.data30(data30),
.data31(data31),
.clk(clk),
.rst_n(rst_n),
.buffer0(buffer0),
.buffer1(buffer1),
.buffer2(buffer2),
.buffer3(buffer3),
.buffer4(buffer4),
.buffer5(buffer5),
.buffer6(buffer6),
.buffer7(buffer7),
.buffer8(buffer8),
.buffer9(buffer9),
.buffer10(buffer10),
.buffer11(buffer11),
.buffer12(buffer12),
.buffer13(buffer13),
.buffer14(buffer14),
.buffer15(buffer15),
.buffer16(buffer16),
.buffer17(buffer17),
.buffer18(buffer18),
.buffer19(buffer19),
.buffer20(buffer20),
.buffer21(buffer21),
.buffer22(buffer22),
.buffer23(buffer23),
.buffer24(buffer24),
.buffer25(buffer25),
.buffer26(buffer26),
.buffer27(buffer27),
.buffer28(buffer28),
.buffer29(buffer29),
.buffer30(buffer30),
.buffer31(buffer31),
.valid_out(valid_out_input_buffer)
);

zero_padding_second #(
.DATA_WIDTH(32),
.PAD_WIDTH(15),
.PAD_HEIGHT(19),
.WIDTH(13),
.HEIGHT(17)
)zero_padding_second(
 .buffer0(buffer0),
.buffer1(buffer1),
.buffer2(buffer2),
.buffer3(buffer3),
.buffer4(buffer4),
.buffer5(buffer5),
.buffer6(buffer6),
.buffer7(buffer7),
.buffer8(buffer8),
.buffer9(buffer9),
.buffer10(buffer10),
.buffer11(buffer11),
.buffer12(buffer12),
.buffer13(buffer13),
.buffer14(buffer14),
.buffer15(buffer15),
.buffer16(buffer16),
.buffer17(buffer17),
.buffer18(buffer18),
.buffer19(buffer19),
.buffer20(buffer20),
.buffer21(buffer21),
.buffer22(buffer22),
.buffer23(buffer23),
.buffer24(buffer24),
.buffer25(buffer25),
.buffer26(buffer26),
.buffer27(buffer27),
.buffer28(buffer28),
.buffer29(buffer29),
.buffer30(buffer30),
.buffer31(buffer31),
.valid_in(valid_out_input_buffer),
.rst_n(rst_n),
.clk(clk),
.padded0(padded0),
.padded1(padded1),
.padded2(padded2),
.padded3(padded3),
.padded4(padded4),
.padded5(padded5),
.padded6(padded6),
.padded7(padded7),
.padded8(padded8),
.padded9(padded9),
.padded10(padded10),
.padded11(padded11),
.padded12(padded12),
.padded13(padded13),
.padded14(padded14),
.padded15(padded15),
.padded16(padded16),
.padded17(padded17),
.padded18(padded18),
.padded19(padded19),
.padded20(padded20),
.padded21(padded21),
.padded22(padded22),
.padded23(padded23),
.padded24(padded24),
.padded25(padded25),
.padded26(padded26),
.padded27(padded27),
.padded28(padded28),
.padded29(padded29),
.padded30(padded30),
.padded31(padded31),
.valid_padding(valid_out_zero_padding_second)
);

threebythree #(
.DATA_WIDTH(32),
.PAD_WIDTH(15),
.PAD_HEIGHT(19)
)threebythree(
.padded0(padded0),
.padded1(padded1),
.padded2(padded2),
.padded3(padded3),
.padded4(padded4),
.padded5(padded5),
.padded6(padded6),
.padded7(padded7),
.padded8(padded8),
.padded9(padded9),
.padded10(padded10),
.padded11(padded11),
.padded12(padded12),
.padded13(padded13),
.padded14(padded14),
.padded15(padded15),
.padded16(padded16),
.padded17(padded17),
.padded18(padded18),
.padded19(padded19),
.padded20(padded20),
.padded21(padded21),
.padded22(padded22),
.padded23(padded23),
.padded24(padded24),
.padded25(padded25),
.padded26(padded26),
.padded27(padded27),
.padded28(padded28),
.padded29(padded29),
.padded30(padded30),
.padded31(padded31),
.valid_padding(valid_out_zero_padding_second),
.rst_n(rst_n),
.clk(clk),
.patch(patch),
.valid_out(valid_out_threebythree)
);

conv2_layer conv2_layer(
.clk(clk),
.rst_n(rst_n),
.valid_in(valid_out_threebythree),
.data_in(patch),
.conv2_out(data_out_conv2),
.valid_out(valid_out_conv2)
);

conv2_accum #(
.WIDTH(13),
.HEIGHT(17),
.SIZE(221),
.filter_num(64),
.channel_num(32)
) conv2_accum(
.data_in(data_out_conv2),
.valid_in(valid_out_conv2),
.clk(clk),
.rst_n(rst_n),
.data_out(data_out_conv2_accum),
.valid_out(valid_out_conv2_accum)
);

relu2#(
.IMAGE_WIDTH(13),
.IMAGE_HEIGHT(17),
.CHANNELS(64),
.DATA_BITS(32)
)relu2(
.data_in(data_out_conv2_accum),
.valid_in(valid_out_conv2_accum),
.rst_n(rst_n),
.clk(clk),
.data_out(data_out_relu2),
.valid_out(valid_out_relu2)
);

channel_buffer2#(
.IMAGE_WIDTH(13),
.IMAGE_HEIGHT(17),
.CHANNELS(64),
.DATA_BITS(32)
)channel_buffer2(
.data_in(data_out_relu2),
.valid_in(valid_out_relu2),
.clk(clk),
.rst_n(rst_n),
.data_out_1(data_out_buf_1),
.data_out_2(data_out_buf_2),
.data_out_3(data_out_buf_3),
.data_out_4(data_out_buf_4),
.data_out_5(data_out_buf_5),
.data_out_6(data_out_buf_6),
.data_out_7(data_out_buf_7),
.data_out_8(data_out_buf_8),
.data_out_9(data_out_buf_9),
.data_out_10(data_out_buf_10),
.data_out_11(data_out_buf_11),
.data_out_12(data_out_buf_12),
.data_out_13(data_out_buf_13),
.data_out_14(data_out_buf_14),
.data_out_15(data_out_buf_15),
.data_out_16(data_out_buf_16),
.data_out_17(data_out_buf_17),
.data_out_18(data_out_buf_18),
.data_out_19(data_out_buf_19),
.data_out_20(data_out_buf_20),
.data_out_21(data_out_buf_21),
.data_out_22(data_out_buf_22),
.data_out_23(data_out_buf_23),
.data_out_24(data_out_buf_24),
.data_out_25(data_out_buf_25),
.data_out_26(data_out_buf_26),
.data_out_27(data_out_buf_27),
.data_out_28(data_out_buf_28),
.data_out_29(data_out_buf_29),
.data_out_30(data_out_buf_30),
.data_out_31(data_out_buf_31),
.data_out_32(data_out_buf_32),
.data_out_33(data_out_buf_33),
.data_out_34(data_out_buf_34),
.data_out_35(data_out_buf_35),
.data_out_36(data_out_buf_36),
.data_out_37(data_out_buf_37),
.data_out_38(data_out_buf_38),
.data_out_39(data_out_buf_39),
.data_out_40(data_out_buf_40),
.data_out_41(data_out_buf_41),
.data_out_42(data_out_buf_42),
.data_out_43(data_out_buf_43),
.data_out_44(data_out_buf_44),
.data_out_45(data_out_buf_45),
.data_out_46(data_out_buf_46),
.data_out_47(data_out_buf_47),
.data_out_48(data_out_buf_48),
.data_out_49(data_out_buf_49),
.data_out_50(data_out_buf_50),
.data_out_51(data_out_buf_51),
.data_out_52(data_out_buf_52),
.data_out_53(data_out_buf_53),
.data_out_54(data_out_buf_54),
.data_out_55(data_out_buf_55),
.data_out_56(data_out_buf_56),
.data_out_57(data_out_buf_57),
.data_out_58(data_out_buf_58),
.data_out_59(data_out_buf_59),
.data_out_60(data_out_buf_60),
.data_out_61(data_out_buf_61),
.data_out_62(data_out_buf_62),
.data_out_63(data_out_buf_63),
.data_out_64(data_out_buf_64),
.valid_out(valid_out_channel_buffer2)
);

max_pooling_layer_top2 max_pooling_layer_top2(
.valid_in(valid_out_channel_buffer2),
.rst_n(rst_n),
.clk(clk),
.valid_out(valid_out_layer2),
.data_in_1(data_out_buf_1),
.data_in_2(data_out_buf_2),
.data_in_3(data_out_buf_3),
.data_in_4(data_out_buf_4),
.data_in_5(data_out_buf_5),
.data_in_6(data_out_buf_6),
.data_in_7(data_out_buf_7),
.data_in_8(data_out_buf_8),
.data_in_9(data_out_buf_9),
.data_in_10(data_out_buf_10),
.data_in_11(data_out_buf_11),
.data_in_12(data_out_buf_12),
.data_in_13(data_out_buf_13),
.data_in_14(data_out_buf_14),
.data_in_15(data_out_buf_15),
.data_in_16(data_out_buf_16),
.data_in_17(data_out_buf_17),
.data_in_18(data_out_buf_18),
.data_in_19(data_out_buf_19),
.data_in_20(data_out_buf_20),
.data_in_21(data_out_buf_21),
.data_in_22(data_out_buf_22),
.data_in_23(data_out_buf_23),
.data_in_24(data_out_buf_24),
.data_in_25(data_out_buf_25),
.data_in_26(data_out_buf_26),
.data_in_27(data_out_buf_27),
.data_in_28(data_out_buf_28),
.data_in_29(data_out_buf_29),
.data_in_30(data_out_buf_30),
.data_in_31(data_out_buf_31),
.data_in_32(data_out_buf_32),
.data_in_33(data_out_buf_33),
.data_in_34(data_out_buf_34),
.data_in_35(data_out_buf_35),
.data_in_36(data_out_buf_36),
.data_in_37(data_out_buf_37),
.data_in_38(data_out_buf_38),
.data_in_39(data_out_buf_39),
.data_in_40(data_out_buf_40),
.data_in_41(data_out_buf_41),
.data_in_42(data_out_buf_42),
.data_in_43(data_out_buf_43),
.data_in_44(data_out_buf_44),
.data_in_45(data_out_buf_45),
.data_in_46(data_out_buf_46),
.data_in_47(data_out_buf_47),
.data_in_48(data_out_buf_48),
.data_in_49(data_out_buf_49),
.data_in_50(data_out_buf_50),
.data_in_51(data_out_buf_51),
.data_in_52(data_out_buf_52),
.data_in_53(data_out_buf_53),
.data_in_54(data_out_buf_54),
.data_in_55(data_out_buf_55),
.data_in_56(data_out_buf_56),
.data_in_57(data_out_buf_57),
.data_in_58(data_out_buf_58),
.data_in_59(data_out_buf_59),
.data_in_60(data_out_buf_60),
.data_in_61(data_out_buf_61),
.data_in_62(data_out_buf_62),
.data_in_63(data_out_buf_63),
.data_in_64(data_out_buf_64),
.data_out_1(data_out_1),
.data_out_2(data_out_2),
.data_out_3(data_out_3),
.data_out_4(data_out_4),
.data_out_5(data_out_5),
.data_out_6(data_out_6),
.data_out_7(data_out_7),
.data_out_8(data_out_8),
.data_out_9(data_out_9),
.data_out_10(data_out_10),
.data_out_11(data_out_11),
.data_out_12(data_out_12),
.data_out_13(data_out_13),
.data_out_14(data_out_14),
.data_out_15(data_out_15),
.data_out_16(data_out_16),
.data_out_17(data_out_17),
.data_out_18(data_out_18),
.data_out_19(data_out_19),
.data_out_20(data_out_20),
.data_out_21(data_out_21),
.data_out_22(data_out_22),
.data_out_23(data_out_23),
.data_out_24(data_out_24),
.data_out_25(data_out_25),
.data_out_26(data_out_26),
.data_out_27(data_out_27),
.data_out_28(data_out_28),
.data_out_29(data_out_29),
.data_out_30(data_out_30),
.data_out_31(data_out_31),
.data_out_32(data_out_32),
.data_out_33(data_out_33),
.data_out_34(data_out_34),
.data_out_35(data_out_35),
.data_out_36(data_out_36),
.data_out_37(data_out_37),
.data_out_38(data_out_38),
.data_out_39(data_out_39),
.data_out_40(data_out_40),
.data_out_41(data_out_41),
.data_out_42(data_out_42),
.data_out_43(data_out_43),
.data_out_44(data_out_44),
.data_out_45(data_out_45),
.data_out_46(data_out_46),
.data_out_47(data_out_47),
.data_out_48(data_out_48),
.data_out_49(data_out_49),
.data_out_50(data_out_50),
.data_out_51(data_out_51),
.data_out_52(data_out_52),
.data_out_53(data_out_53),
.data_out_54(data_out_54),
.data_out_55(data_out_55),
.data_out_56(data_out_56),
.data_out_57(data_out_57),
.data_out_58(data_out_58),
.data_out_59(data_out_59),
.data_out_60(data_out_60),
.data_out_61(data_out_61),
.data_out_62(data_out_62),
.data_out_63(data_out_63),
.data_out_64(data_out_64)
);

endmodule
